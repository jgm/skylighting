architecture arch of device is
begin
    process
    begin
    end process;
end arch;
